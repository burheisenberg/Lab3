----------------------------------------------------------------------------------
-- COMPANY: 	KOC UNIVERSITY
-- ENGINEER: 	ONURHAN OZTURK
-- 
-- CREATE DATE:    18:21:21 04/26/2016 
-- DESIGN NAME: 	
-- MODULE NAME:    SEVSEG_DECODER - BEHAVIORAL 
-- PROJECT NAME: 	 SSSLIB
-- TARGET DEVICES: SPARTAN 3E
-- TOOL VERSIONS: 
-- DESCRIPTION: 
--
-- DEPENDENCIES: 
--
-- REVISION: 
-- REVISION 0.01 - FILE CREATED
-- ADDITIONAL COMMENTS: 
--
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- UNCOMMENT THE FOLLOWING LIBRARY DECLARATION IF USING
-- ARITHMETIC FUNCTIONS WITH SIGNED OR UNSIGNED VALUES
--USE IEEE.NUMERIC_STD.ALL;

-- UNCOMMENT THE FOLLOWING LIBRARY DECLARATION IF INSTANTIATING
-- ANY XILINX PRIMITIVES IN THIS CODE.
--LIBRARY UNISIM;
--USE UNISIM.VCOMPONENTS.ALL;

ENTITY SEVSEG_DECODER IS
    PORT ( INPUT : IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
           SEVSEG_BUS : OUT  STD_LOGIC_VECTOR (6 DOWNTO 0));
END SEVSEG_DECODER;

ARCHITECTURE BEHAVIORAL OF SEVSEG_DECODER IS

BEGIN

WITH INPUT SELECT SEVSEG_BUS <=
	"0000001" WHEN "0000", --0
	"1001111" WHEN "0001", --1
	"0010010" WHEN "0010", --2
	"0000110" WHEN "0011", --3
	"1001100" WHEN "0100", --4
	"0100100" WHEN "0101", --5
	"0100000" WHEN "0110", --6
	"0001111" WHEN "0111", --7
	"0000000" WHEN "1000", --8
	"0001111" WHEN "1001", --7
	"0100000" WHEN "1010", --6
	"0100100" WHEN "1011", --5
	"1001100" WHEN "1100", --4
	"0000110" WHEN "1101", --3
	"0010010" WHEN "1110", --2
	"1001111" WHEN "1111", --1
	"0000001" WHEN OTHERS;
END BEHAVIORAL;

